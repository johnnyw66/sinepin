// SineROM case statement was generated using a simple
// bit of python. This table is a quarter of a sine wave.

/*

import math ;

fpmult <= 32768 ;		#16bit
for i in range (256):
    a <= i ;	
    sv <= ( 1 +  math.sin(a * math.pi / 512)) ;
    fpsv <=  int(fpmult * sv) ;
    # print("%d %d %d" % (i,fpsv, int(fpsv / 256))) ;
    print("8'd%d : svalue <= 16'd%d ;" % (i,fpsv)) ;

*/

module sineQuartROM #(parameter SINEROMSIZE = 1024)(
	input clk,
	input [7:0] address,
	output reg [15:0] svalue
);


always @(posedge clk)
begin
	case(address)
		8'd0 : svalue <= 16'd32768 ;
		8'd1 : svalue <= 16'd32969 ;
		8'd2 : svalue <= 16'd33170 ;
		8'd3 : svalue <= 16'd33371 ;
		8'd4 : svalue <= 16'd33572 ;
		8'd5 : svalue <= 16'd33773 ;
		8'd6 : svalue <= 16'd33974 ;
		8'd7 : svalue <= 16'd34175 ;
		8'd8 : svalue <= 16'd34375 ;
		8'd9 : svalue <= 16'd34576 ;
		8'd10 : svalue <= 16'd34777 ;
		8'd11 : svalue <= 16'd34978 ;
		8'd12 : svalue <= 16'd35178 ;
		8'd13 : svalue <= 16'd35379 ;
		8'd14 : svalue <= 16'd35579 ;
		8'd15 : svalue <= 16'd35779 ;
		8'd16 : svalue <= 16'd35979 ;
		8'd17 : svalue <= 16'd36179 ;
		8'd18 : svalue <= 16'd36379 ;
		8'd19 : svalue <= 16'd36579 ;
		8'd20 : svalue <= 16'd36779 ;
		8'd21 : svalue <= 16'd36978 ;
		8'd22 : svalue <= 16'd37177 ;
		8'd23 : svalue <= 16'd37377 ;
		8'd24 : svalue <= 16'd37576 ;
		8'd25 : svalue <= 16'd37774 ;
		8'd26 : svalue <= 16'd37973 ;
		8'd27 : svalue <= 16'd38171 ;
		8'd28 : svalue <= 16'd38370 ;
		8'd29 : svalue <= 16'd38568 ;
		8'd30 : svalue <= 16'd38765 ;
		8'd31 : svalue <= 16'd38963 ;
		8'd32 : svalue <= 16'd39160 ;
		8'd33 : svalue <= 16'd39357 ;
		8'd34 : svalue <= 16'd39554 ;
		8'd35 : svalue <= 16'd39751 ;
		8'd36 : svalue <= 16'd39947 ;
		8'd37 : svalue <= 16'd40143 ;
		8'd38 : svalue <= 16'd40339 ;
		8'd39 : svalue <= 16'd40534 ;
		8'd40 : svalue <= 16'd40729 ;
		8'd41 : svalue <= 16'd40924 ;
		8'd42 : svalue <= 16'd41119 ;
		8'd43 : svalue <= 16'd41313 ;
		8'd44 : svalue <= 16'd41507 ;
		8'd45 : svalue <= 16'd41701 ;
		8'd46 : svalue <= 16'd41894 ;
		8'd47 : svalue <= 16'd42087 ;
		8'd48 : svalue <= 16'd42280 ;
		8'd49 : svalue <= 16'd42472 ;
		8'd50 : svalue <= 16'd42664 ;
		8'd51 : svalue <= 16'd42855 ;
		8'd52 : svalue <= 16'd43046 ;
		8'd53 : svalue <= 16'd43237 ;
		8'd54 : svalue <= 16'd43427 ;
		8'd55 : svalue <= 16'd43617 ;
		8'd56 : svalue <= 16'd43807 ;
		8'd57 : svalue <= 16'd43996 ;
		8'd58 : svalue <= 16'd44184 ;
		8'd59 : svalue <= 16'd44373 ;
		8'd60 : svalue <= 16'd44561 ;
		8'd61 : svalue <= 16'd44748 ;
		8'd62 : svalue <= 16'd44935 ;
		8'd63 : svalue <= 16'd45121 ;
		8'd64 : svalue <= 16'd45307 ;
		8'd65 : svalue <= 16'd45493 ;
		8'd66 : svalue <= 16'd45678 ;
		8'd67 : svalue <= 16'd45862 ;
		8'd68 : svalue <= 16'd46046 ;
		8'd69 : svalue <= 16'd46230 ;
		8'd70 : svalue <= 16'd46413 ;
		8'd71 : svalue <= 16'd46596 ;
		8'd72 : svalue <= 16'd46778 ;
		8'd73 : svalue <= 16'd46959 ;
		8'd74 : svalue <= 16'd47140 ;
		8'd75 : svalue <= 16'd47320 ;
		8'd76 : svalue <= 16'd47500 ;
		8'd77 : svalue <= 16'd47680 ;
		8'd78 : svalue <= 16'd47858 ;
		8'd79 : svalue <= 16'd48037 ;
		8'd80 : svalue <= 16'd48214 ;
		8'd81 : svalue <= 16'd48391 ;
		8'd82 : svalue <= 16'd48568 ;
		8'd83 : svalue <= 16'd48744 ;
		8'd84 : svalue <= 16'd48919 ;
		8'd85 : svalue <= 16'd49093 ;
		8'd86 : svalue <= 16'd49267 ;
		8'd87 : svalue <= 16'd49441 ;
		8'd88 : svalue <= 16'd49614 ;
		8'd89 : svalue <= 16'd49786 ;
		8'd90 : svalue <= 16'd49957 ;
		8'd91 : svalue <= 16'd50128 ;
		8'd92 : svalue <= 16'd50298 ;
		8'd93 : svalue <= 16'd50468 ;
		8'd94 : svalue <= 16'd50637 ;
		8'd95 : svalue <= 16'd50805 ;
		8'd96 : svalue <= 16'd50972 ;
		8'd97 : svalue <= 16'd51139 ;
		8'd98 : svalue <= 16'd51305 ;
		8'd99 : svalue <= 16'd51471 ;
		8'd100 : svalue <= 16'd51636 ;
		8'd101 : svalue <= 16'd51800 ;
		8'd102 : svalue <= 16'd51963 ;
		8'd103 : svalue <= 16'd52126 ;
		8'd104 : svalue <= 16'd52287 ;
		8'd105 : svalue <= 16'd52449 ;
		8'd106 : svalue <= 16'd52609 ;
		8'd107 : svalue <= 16'd52769 ;
		8'd108 : svalue <= 16'd52927 ;
		8'd109 : svalue <= 16'd53086 ;
		8'd110 : svalue <= 16'd53243 ;
		8'd111 : svalue <= 16'd53399 ;
		8'd112 : svalue <= 16'd53555 ;
		8'd113 : svalue <= 16'd53710 ;
		8'd114 : svalue <= 16'd53865 ;
		8'd115 : svalue <= 16'd54018 ;
		8'd116 : svalue <= 16'd54171 ;
		8'd117 : svalue <= 16'd54323 ;
		8'd118 : svalue <= 16'd54474 ;
		8'd119 : svalue <= 16'd54624 ;
		8'd120 : svalue <= 16'd54773 ;
		8'd121 : svalue <= 16'd54922 ;
		8'd122 : svalue <= 16'd55069 ;
		8'd123 : svalue <= 16'd55216 ;
		8'd124 : svalue <= 16'd55362 ;
		8'd125 : svalue <= 16'd55508 ;
		8'd126 : svalue <= 16'd55652 ;
		8'd127 : svalue <= 16'd55795 ;
		8'd128 : svalue <= 16'd55938 ;
		8'd129 : svalue <= 16'd56080 ;
		8'd130 : svalue <= 16'd56221 ;
		8'd131 : svalue <= 16'd56361 ;
		8'd132 : svalue <= 16'd56500 ;
		8'd133 : svalue <= 16'd56638 ;
		8'd134 : svalue <= 16'd56775 ;
		8'd135 : svalue <= 16'd56912 ;
		8'd136 : svalue <= 16'd57047 ;
		8'd137 : svalue <= 16'd57182 ;
		8'd138 : svalue <= 16'd57315 ;
		8'd139 : svalue <= 16'd57448 ;
		8'd140 : svalue <= 16'd57580 ;
		8'd141 : svalue <= 16'd57711 ;
		8'd142 : svalue <= 16'd57841 ;
		8'd143 : svalue <= 16'd57969 ;
		8'd144 : svalue <= 16'd58098 ;
		8'd145 : svalue <= 16'd58225 ;
		8'd146 : svalue <= 16'd58351 ;
		8'd147 : svalue <= 16'd58476 ;
		8'd148 : svalue <= 16'd58600 ;
		8'd149 : svalue <= 16'd58723 ;
		8'd150 : svalue <= 16'd58845 ;
		8'd151 : svalue <= 16'd58967 ;
		8'd152 : svalue <= 16'd59087 ;
		8'd153 : svalue <= 16'd59206 ;
		8'd154 : svalue <= 16'd59325 ;
		8'd155 : svalue <= 16'd59442 ;
		8'd156 : svalue <= 16'd59558 ;
		8'd157 : svalue <= 16'd59673 ;
		8'd158 : svalue <= 16'd59788 ;
		8'd159 : svalue <= 16'd59901 ;
		8'd160 : svalue <= 16'd60013 ;
		8'd161 : svalue <= 16'd60124 ;
		8'd162 : svalue <= 16'd60234 ;
		8'd163 : svalue <= 16'd60344 ;
		8'd164 : svalue <= 16'd60452 ;
		8'd165 : svalue <= 16'd60559 ;
		8'd166 : svalue <= 16'd60665 ;
		8'd167 : svalue <= 16'd60770 ;
		8'd168 : svalue <= 16'd60874 ;
		8'd169 : svalue <= 16'd60976 ;
		8'd170 : svalue <= 16'd61078 ;
		8'd171 : svalue <= 16'd61179 ;
		8'd172 : svalue <= 16'd61279 ;
		8'd173 : svalue <= 16'd61377 ;
		8'd174 : svalue <= 16'd61475 ;
		8'd175 : svalue <= 16'd61571 ;
		8'd176 : svalue <= 16'd61666 ;
		8'd177 : svalue <= 16'd61761 ;
		8'd178 : svalue <= 16'd61854 ;
		8'd179 : svalue <= 16'd61946 ;
		8'd180 : svalue <= 16'd62037 ;
		8'd181 : svalue <= 16'd62127 ;
		8'd182 : svalue <= 16'd62215 ;
		8'd183 : svalue <= 16'd62303 ;
		8'd184 : svalue <= 16'd62389 ;
		8'd185 : svalue <= 16'd62475 ;
		8'd186 : svalue <= 16'd62559 ;
		8'd187 : svalue <= 16'd62642 ;
		8'd188 : svalue <= 16'd62724 ;
		8'd189 : svalue <= 16'd62805 ;
		8'd190 : svalue <= 16'd62885 ;
		8'd191 : svalue <= 16'd62964 ;
		8'd192 : svalue <= 16'd63041 ;
		8'd193 : svalue <= 16'd63118 ;
		8'd194 : svalue <= 16'd63193 ;
		8'd195 : svalue <= 16'd63267 ;
		8'd196 : svalue <= 16'd63340 ;
		8'd197 : svalue <= 16'd63412 ;
		8'd198 : svalue <= 16'd63482 ;
		8'd199 : svalue <= 16'd63552 ;
		8'd200 : svalue <= 16'd63620 ;
		8'd201 : svalue <= 16'd63687 ;
		8'd202 : svalue <= 16'd63753 ;
		8'd203 : svalue <= 16'd63818 ;
		8'd204 : svalue <= 16'd63882 ;
		8'd205 : svalue <= 16'd63944 ;
		8'd206 : svalue <= 16'd64005 ;
		8'd207 : svalue <= 16'd64066 ;
		8'd208 : svalue <= 16'd64125 ;
		8'd209 : svalue <= 16'd64182 ;
		8'd210 : svalue <= 16'd64239 ;
		8'd211 : svalue <= 16'd64294 ;
		8'd212 : svalue <= 16'd64349 ;
		8'd213 : svalue <= 16'd64402 ;
		8'd214 : svalue <= 16'd64453 ;
		8'd215 : svalue <= 16'd64504 ;
		8'd216 : svalue <= 16'd64553 ;
		8'd217 : svalue <= 16'd64602 ;
		8'd218 : svalue <= 16'd64649 ;
		8'd219 : svalue <= 16'd64695 ;
		8'd220 : svalue <= 16'd64739 ;
		8'd221 : svalue <= 16'd64783 ;
		8'd222 : svalue <= 16'd64825 ;
		8'd223 : svalue <= 16'd64866 ;
		8'd224 : svalue <= 16'd64906 ;
		8'd225 : svalue <= 16'd64944 ;
		8'd226 : svalue <= 16'd64982 ;
		8'd227 : svalue <= 16'd65018 ;
		8'd228 : svalue <= 16'd65053 ;
		8'd229 : svalue <= 16'd65087 ;
		8'd230 : svalue <= 16'd65119 ;
		8'd231 : svalue <= 16'd65151 ;
		8'd232 : svalue <= 16'd65181 ;
		8'd233 : svalue <= 16'd65210 ;
		8'd234 : svalue <= 16'd65237 ;
		8'd235 : svalue <= 16'd65264 ;
		8'd236 : svalue <= 16'd65289 ;
		8'd237 : svalue <= 16'd65313 ;
		8'd238 : svalue <= 16'd65336 ;
		8'd239 : svalue <= 16'd65357 ;
		8'd240 : svalue <= 16'd65378 ;
		8'd241 : svalue <= 16'd65397 ;
		8'd242 : svalue <= 16'd65415 ;
		8'd243 : svalue <= 16'd65431 ;
		8'd244 : svalue <= 16'd65447 ;
		8'd245 : svalue <= 16'd65461 ;
		8'd246 : svalue <= 16'd65474 ;
		8'd247 : svalue <= 16'd65486 ;
		8'd248 : svalue <= 16'd65496 ;
		8'd249 : svalue <= 16'd65505 ;
		8'd250 : svalue <= 16'd65513 ;
		8'd251 : svalue <= 16'd65520 ;
		8'd252 : svalue <= 16'd65526 ;
		8'd253 : svalue <= 16'd65530 ;
		8'd254 : svalue <= 16'd65533 ;
		8'd255 : svalue <= 16'd65535 ;
			
	endcase
	
end

endmodule
