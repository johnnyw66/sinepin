module musicMarioROM2  (
	input clk,
	input [8:0] address,
	output reg [7:0] note
);

always @(posedge clk)
	
	case(address[8:0])
			0: note <= 8'd66 ;
			1: note <= 8'd66 ;
			2: note <= 8'd255 ;
			3: note <= 8'd66 ;
			4: note <= 8'd255 ;
			5: note <= 8'd66 ;
			6: note <= 8'd66 ;
			7: note <= 8'd255 ;
			8: note <= 8'd71 ;
			9: note <= 8'd255 ;
			10: note <= 8'd255 ;
			11: note <= 8'd255 ;
			12: note <= 8'd67 ;
			13: note <= 8'd255 ;
			14: note <= 8'd255 ;
			15: note <= 8'd255 ;
			16: note <= 8'd64 ;
			17: note <= 8'd255 ;
			18: note <= 8'd255 ;
			19: note <= 8'd60 ;
			20: note <= 8'd255 ;
			21: note <= 8'd255 ;
			22: note <= 8'd55 ;
			23: note <= 8'd255 ;
			24: note <= 8'd255 ;
			25: note <= 8'd60 ;
			26: note <= 8'd255 ;
			27: note <= 8'd62 ;
			28: note <= 8'd255 ;
			29: note <= 8'd61 ;
			30: note <= 8'd60 ;
			31: note <= 8'd255 ;
			32: note <= 8'd60 ;
			33: note <= 8'd67 ;
			34: note <= 8'd71 ;
			35: note <= 8'd72 ;
			36: note <= 8'd255 ;
			37: note <= 8'd69 ;
			38: note <= 8'd71 ;
			39: note <= 8'd255 ;
			40: note <= 8'd69 ;
			41: note <= 8'd255 ;
			42: note <= 8'd64 ;
			43: note <= 8'd65 ;
			44: note <= 8'd62 ;
			45: note <= 8'd255 ;
			46: note <= 8'd255 ;
			47: note <= 8'd64 ;
			48: note <= 8'd255 ;
			49: note <= 8'd255 ;
			50: note <= 8'd60 ;
			51: note <= 8'd255 ;
			52: note <= 8'd255 ;
			53: note <= 8'd55 ;
			54: note <= 8'd255 ;
			55: note <= 8'd255 ;
			56: note <= 8'd60 ;
			57: note <= 8'd255 ;
			58: note <= 8'd62 ;
			59: note <= 8'd255 ;
			60: note <= 8'd61 ;
			61: note <= 8'd60 ;
			62: note <= 8'd255 ;
			63: note <= 8'd60 ;
			64: note <= 8'd67 ;
			65: note <= 8'd71 ;
			66: note <= 8'd72 ;
			67: note <= 8'd255 ;
			68: note <= 8'd69 ;
			69: note <= 8'd71 ;
			70: note <= 8'd255 ;
			71: note <= 8'd69 ;
			72: note <= 8'd255 ;
			73: note <= 8'd64 ;
			74: note <= 8'd65 ;
			75: note <= 8'd62 ;
			76: note <= 8'd255 ;
			77: note <= 8'd255 ;
			78: note <= 8'd255 ;
			79: note <= 8'd255 ;
			80: note <= 8'd76 ;
			81: note <= 8'd75 ;
			82: note <= 8'd74 ;
			83: note <= 8'd71 ;
			84: note <= 8'd255 ;
			85: note <= 8'd72 ;
			86: note <= 8'd255 ;
			87: note <= 8'd64 ;
			88: note <= 8'd65 ;
			89: note <= 8'd67 ;
			90: note <= 8'd255 ;
			91: note <= 8'd60 ;
			92: note <= 8'd64 ;
			93: note <= 8'd65 ;
			94: note <= 8'd255 ;
			95: note <= 8'd255 ;
			96: note <= 8'd76 ;
			97: note <= 8'd75 ;
			98: note <= 8'd74 ;
			99: note <= 8'd71 ;
			100: note <= 8'd255 ;
			101: note <= 8'd72 ;
			102: note <= 8'd255 ;
			103: note <= 8'd77 ;
			104: note <= 8'd255 ;
			105: note <= 8'd77 ;
			106: note <= 8'd77 ;
			107: note <= 8'd255 ;
			108: note <= 8'd255 ;
			109: note <= 8'd255 ;
			110: note <= 8'd255 ;
			111: note <= 8'd255 ;
			112: note <= 8'd76 ;
			113: note <= 8'd75 ;
			114: note <= 8'd74 ;
			115: note <= 8'd71 ;
			116: note <= 8'd255 ;
			117: note <= 8'd72 ;
			118: note <= 8'd255 ;
			119: note <= 8'd64 ;
			120: note <= 8'd65 ;
			121: note <= 8'd67 ;
			122: note <= 8'd255 ;
			123: note <= 8'd60 ;
			124: note <= 8'd64 ;
			125: note <= 8'd65 ;
			126: note <= 8'd255 ;
			127: note <= 8'd255 ;
			128: note <= 8'd68 ;
			129: note <= 8'd255 ;
			130: note <= 8'd255 ;
			131: note <= 8'd65 ;
			132: note <= 8'd255 ;
			133: note <= 8'd255 ;
			134: note <= 8'd64 ;
			135: note <= 8'd255 ;
			136: note <= 8'd255 ;
			137: note <= 8'd255 ;
			138: note <= 8'd255 ;
			139: note <= 8'd255 ;
			140: note <= 8'd255 ;
			141: note <= 8'd255 ;
			142: note <= 8'd255 ;
			143: note <= 8'd255 ;
			144: note <= 8'd76 ;
			145: note <= 8'd75 ;
			146: note <= 8'd74 ;
			147: note <= 8'd71 ;
			148: note <= 8'd255 ;
			149: note <= 8'd72 ;
			150: note <= 8'd255 ;
			151: note <= 8'd64 ;
			152: note <= 8'd65 ;
			153: note <= 8'd67 ;
			154: note <= 8'd255 ;
			155: note <= 8'd60 ;
			156: note <= 8'd64 ;
			157: note <= 8'd65 ;
			158: note <= 8'd255 ;
			159: note <= 8'd255 ;
			160: note <= 8'd76 ;
			161: note <= 8'd75 ;
			162: note <= 8'd74 ;
			163: note <= 8'd71 ;
			164: note <= 8'd255 ;
			165: note <= 8'd72 ;
			166: note <= 8'd255 ;
			167: note <= 8'd77 ;
			168: note <= 8'd255 ;
			169: note <= 8'd77 ;
			170: note <= 8'd77 ;
			171: note <= 8'd255 ;
			172: note <= 8'd255 ;
			173: note <= 8'd255 ;
			174: note <= 8'd255 ;
			175: note <= 8'd255 ;
			176: note <= 8'd76 ;
			177: note <= 8'd75 ;
			178: note <= 8'd74 ;
			179: note <= 8'd71 ;
			180: note <= 8'd255 ;
			181: note <= 8'd72 ;
			182: note <= 8'd255 ;
			183: note <= 8'd64 ;
			184: note <= 8'd65 ;
			185: note <= 8'd67 ;
			186: note <= 8'd255 ;
			187: note <= 8'd60 ;
			188: note <= 8'd64 ;
			189: note <= 8'd65 ;
			190: note <= 8'd255 ;
			191: note <= 8'd255 ;
			192: note <= 8'd68 ;
			193: note <= 8'd255 ;
			194: note <= 8'd255 ;
			195: note <= 8'd65 ;
			196: note <= 8'd255 ;
			197: note <= 8'd255 ;
			198: note <= 8'd64 ;
			199: note <= 8'd255 ;
			200: note <= 8'd255 ;
			201: note <= 8'd255 ;
			202: note <= 8'd255 ;
			203: note <= 8'd255 ;
			204: note <= 8'd255 ;
			205: note <= 8'd255 ;
			206: note <= 8'd68 ;
			207: note <= 8'd68 ;
			208: note <= 8'd255 ;
			209: note <= 8'd68 ;
			210: note <= 8'd255 ;
			211: note <= 8'd68 ;
			212: note <= 8'd70 ;
			213: note <= 8'd255 ;
			214: note <= 8'd67 ;
			215: note <= 8'd64 ;
			216: note <= 8'd255 ;
			217: note <= 8'd64 ;
			218: note <= 8'd60 ;
			219: note <= 8'd255 ;
			220: note <= 8'd255 ;
			221: note <= 8'd255 ;
			222: note <= 8'd68 ;
			223: note <= 8'd68 ;
			224: note <= 8'd255 ;
			225: note <= 8'd68 ;
			226: note <= 8'd255 ;
			227: note <= 8'd68 ;
			228: note <= 8'd70 ;
			229: note <= 8'd67 ;
			230: note <= 8'd255 ;
			231: note <= 8'd255 ;
			232: note <= 8'd255 ;
			233: note <= 8'd255 ;
			234: note <= 8'd255 ;
			235: note <= 8'd255 ;
			236: note <= 8'd255 ;
			237: note <= 8'd255 ;
			238: note <= 8'd68 ;
			239: note <= 8'd68 ;
			240: note <= 8'd255 ;
			241: note <= 8'd68 ;
			242: note <= 8'd255 ;
			243: note <= 8'd68 ;
			244: note <= 8'd70 ;
			245: note <= 8'd255 ;
			246: note <= 8'd67 ;
			247: note <= 8'd64 ;
			248: note <= 8'd255 ;
			249: note <= 8'd64 ;
			250: note <= 8'd60 ;
			251: note <= 8'd255 ;
			252: note <= 8'd255 ;
			253: note <= 8'd255 ;
			254: note <= 8'd66 ;
			255: note <= 8'd66 ;
			256: note <= 8'd255 ;
			257: note <= 8'd66 ;
			258: note <= 8'd255 ;
			259: note <= 8'd66 ;
			260: note <= 8'd66 ;
			261: note <= 8'd255 ;
			262: note <= 8'd71 ;
			263: note <= 8'd255 ;
			264: note <= 8'd255 ;
			265: note <= 8'd255 ;
			266: note <= 8'd67 ;
			267: note <= 8'd255 ;
			268: note <= 8'd255 ;
			269: note <= 8'd255 ;
			270: note <= 8'd72 ;
			271: note <= 8'd69 ;
			272: note <= 8'd255 ;
			273: note <= 8'd64 ;
			274: note <= 8'd255 ;
			275: note <= 8'd255 ;
			276: note <= 8'd64 ;
			277: note <= 8'd255 ;
			278: note <= 8'd65 ;
			279: note <= 8'd72 ;
			280: note <= 8'd255 ;
			281: note <= 8'd72 ;
			282: note <= 8'd65 ;
			283: note <= 8'd255 ;
			284: note <= 8'd255 ;
			285: note <= 8'd255 ;
			286: note <= 8'd67 ;
			287: note <= 8'd77 ;
			288: note <= 8'd77 ;
			289: note <= 8'd77 ;
			290: note <= 8'd76 ;
			291: note <= 8'd74 ;
			292: note <= 8'd72 ;
			293: note <= 8'd69 ;
			294: note <= 8'd255 ;
			295: note <= 8'd65 ;
			296: note <= 8'd64 ;
			297: note <= 8'd255 ;
			298: note <= 8'd255 ;
			299: note <= 8'd255 ;
			300: note <= 8'd72 ;
			301: note <= 8'd69 ;
			302: note <= 8'd255 ;
			303: note <= 8'd64 ;
			304: note <= 8'd255 ;
			305: note <= 8'd255 ;
			306: note <= 8'd64 ;
			307: note <= 8'd255 ;
			308: note <= 8'd65 ;
			309: note <= 8'd72 ;
			310: note <= 8'd255 ;
			311: note <= 8'd72 ;
			312: note <= 8'd65 ;
			313: note <= 8'd255 ;
			314: note <= 8'd255 ;
			315: note <= 8'd255 ;
			316: note <= 8'd67 ;
			317: note <= 8'd74 ;
			318: note <= 8'd255 ;
			319: note <= 8'd74 ;
			320: note <= 8'd74 ;
			321: note <= 8'd72 ;
			322: note <= 8'd71 ;
			323: note <= 8'd72 ;
			324: note <= 8'd255 ;
			325: note <= 8'd255 ;
			326: note <= 8'd255 ;
			327: note <= 8'd255 ;
			328: note <= 8'd255 ;
			329: note <= 8'd255 ;
			330: note <= 8'd255 ;
			default: note <= 8'd1;
	endcase
endmodule
