module powerROM (
	input clk,
	input [7:0] address,
	output  reg [15:0] sinpow
);


always @(posedge clk)
begin
	case(address)
		8'd0 : sinpow <= 0 ;
		8'd1 : sinpow <= 3 ;
		8'd2 : sinpow <= 6 ;
		8'd3 : sinpow <= 8 ;
		8'd4 : sinpow <= 11 ;
		8'd5 : sinpow <= 14 ;
		8'd6 : sinpow <= 17 ;
		8'd7 : sinpow <= 20 ;
		8'd8 : sinpow <= 22 ;
		8'd9 : sinpow <= 25 ;
		8'd10 : sinpow <= 28 ;
		8'd11 : sinpow <= 31 ;
		8'd12 : sinpow <= 34 ;
		8'd13 : sinpow <= 37 ;
		8'd14 : sinpow <= 40 ;
		8'd15 : sinpow <= 42 ;
		8'd16 : sinpow <= 45 ;
		8'd17 : sinpow <= 48 ;
		8'd18 : sinpow <= 51 ;
		8'd19 : sinpow <= 54 ;
		8'd20 : sinpow <= 57 ;
		8'd21 : sinpow <= 60 ;
		8'd22 : sinpow <= 63 ;
		8'd23 : sinpow <= 66 ;
		8'd24 : sinpow <= 69 ;
		8'd25 : sinpow <= 72 ;
		8'd26 : sinpow <= 75 ;
		8'd27 : sinpow <= 78 ;
		8'd28 : sinpow <= 81 ;
		8'd29 : sinpow <= 84 ;
		8'd30 : sinpow <= 87 ;
		8'd31 : sinpow <= 90 ;
		8'd32 : sinpow <= 93 ;
		8'd33 : sinpow <= 96 ;
		8'd34 : sinpow <= 99 ;
		8'd35 : sinpow <= 102 ;
		8'd36 : sinpow <= 105 ;
		8'd37 : sinpow <= 108 ;
		8'd38 : sinpow <= 111 ;
		8'd39 : sinpow <= 114 ;
		8'd40 : sinpow <= 117 ;
		8'd41 : sinpow <= 120 ;
		8'd42 : sinpow <= 123 ;
		8'd43 : sinpow <= 126 ;
		8'd44 : sinpow <= 130 ;
		8'd45 : sinpow <= 133 ;
		8'd46 : sinpow <= 136 ;
		8'd47 : sinpow <= 139 ;
		8'd48 : sinpow <= 142 ;
		8'd49 : sinpow <= 145 ;
		8'd50 : sinpow <= 148 ;
		8'd51 : sinpow <= 152 ;
		8'd52 : sinpow <= 155 ;
		8'd53 : sinpow <= 158 ;
		8'd54 : sinpow <= 161 ;
		8'd55 : sinpow <= 164 ;
		8'd56 : sinpow <= 168 ;
		8'd57 : sinpow <= 171 ;
		8'd58 : sinpow <= 174 ;
		8'd59 : sinpow <= 177 ;
		8'd60 : sinpow <= 181 ;
		8'd61 : sinpow <= 184 ;
		8'd62 : sinpow <= 187 ;
		8'd63 : sinpow <= 190 ;
		8'd64 : sinpow <= 194 ;
		8'd65 : sinpow <= 197 ;
		8'd66 : sinpow <= 200 ;
		8'd67 : sinpow <= 204 ;
		8'd68 : sinpow <= 207 ;
		8'd69 : sinpow <= 210 ;
		8'd70 : sinpow <= 214 ;
		8'd71 : sinpow <= 217 ;
		8'd72 : sinpow <= 220 ;
		8'd73 : sinpow <= 224 ;
		8'd74 : sinpow <= 227 ;
		8'd75 : sinpow <= 231 ;
		8'd76 : sinpow <= 234 ;
		8'd77 : sinpow <= 237 ;
		8'd78 : sinpow <= 241 ;
		8'd79 : sinpow <= 244 ;
		8'd80 : sinpow <= 248 ;
		8'd81 : sinpow <= 251 ;
		8'd82 : sinpow <= 255 ;
		8'd83 : sinpow <= 258 ;
		8'd84 : sinpow <= 262 ;
		8'd85 : sinpow <= 265 ;
		8'd86 : sinpow <= 268 ;
		8'd87 : sinpow <= 272 ;
		8'd88 : sinpow <= 276 ;
		8'd89 : sinpow <= 279 ;
		8'd90 : sinpow <= 283 ;
		8'd91 : sinpow <= 286 ;
		8'd92 : sinpow <= 290 ;
		8'd93 : sinpow <= 293 ;
		8'd94 : sinpow <= 297 ;
		8'd95 : sinpow <= 300 ;
		8'd96 : sinpow <= 304 ;
		8'd97 : sinpow <= 308 ;
		8'd98 : sinpow <= 311 ;
		8'd99 : sinpow <= 315 ;
		8'd100 : sinpow <= 318 ;
		8'd101 : sinpow <= 322 ;
		8'd102 : sinpow <= 326 ;
		8'd103 : sinpow <= 329 ;
		8'd104 : sinpow <= 333 ;
		8'd105 : sinpow <= 337 ;
		8'd106 : sinpow <= 340 ;
		8'd107 : sinpow <= 344 ;
		8'd108 : sinpow <= 348 ;
		8'd109 : sinpow <= 352 ;
		8'd110 : sinpow <= 355 ;
		8'd111 : sinpow <= 359 ;
		8'd112 : sinpow <= 363 ;
		8'd113 : sinpow <= 367 ;
		8'd114 : sinpow <= 370 ;
		8'd115 : sinpow <= 374 ;
		8'd116 : sinpow <= 378 ;
		8'd117 : sinpow <= 382 ;
		8'd118 : sinpow <= 385 ;
		8'd119 : sinpow <= 389 ;
		8'd120 : sinpow <= 393 ;
		8'd121 : sinpow <= 397 ;
		8'd122 : sinpow <= 401 ;
		8'd123 : sinpow <= 405 ;
		8'd124 : sinpow <= 409 ;
		8'd125 : sinpow <= 412 ;
		8'd126 : sinpow <= 416 ;
		8'd127 : sinpow <= 420 ;
		8'd128 : sinpow <= 424 ;
		8'd129 : sinpow <= 428 ;
		8'd130 : sinpow <= 432 ;
		8'd131 : sinpow <= 436 ;
		8'd132 : sinpow <= 440 ;
		8'd133 : sinpow <= 444 ;
		8'd134 : sinpow <= 448 ;
		8'd135 : sinpow <= 452 ;
		8'd136 : sinpow <= 456 ;
		8'd137 : sinpow <= 460 ;
		8'd138 : sinpow <= 464 ;
		8'd139 : sinpow <= 468 ;
		8'd140 : sinpow <= 472 ;
		8'd141 : sinpow <= 476 ;
		8'd142 : sinpow <= 480 ;
		8'd143 : sinpow <= 484 ;
		8'd144 : sinpow <= 488 ;
		8'd145 : sinpow <= 492 ;
		8'd146 : sinpow <= 496 ;
		8'd147 : sinpow <= 501 ;
		8'd148 : sinpow <= 505 ;
		8'd149 : sinpow <= 509 ;
		8'd150 : sinpow <= 513 ;
		8'd151 : sinpow <= 517 ;
		8'd152 : sinpow <= 521 ;
		8'd153 : sinpow <= 526 ;
		8'd154 : sinpow <= 530 ;
		8'd155 : sinpow <= 534 ;
		8'd156 : sinpow <= 538 ;
		8'd157 : sinpow <= 542 ;
		8'd158 : sinpow <= 547 ;
		8'd159 : sinpow <= 551 ;
		8'd160 : sinpow <= 555 ;
		8'd161 : sinpow <= 560 ;
		8'd162 : sinpow <= 564 ;
		8'd163 : sinpow <= 568 ;
		8'd164 : sinpow <= 572 ;
		8'd165 : sinpow <= 577 ;
		8'd166 : sinpow <= 581 ;
		8'd167 : sinpow <= 585 ;
		8'd168 : sinpow <= 590 ;
		8'd169 : sinpow <= 594 ;
		8'd170 : sinpow <= 599 ;
		8'd171 : sinpow <= 603 ;
		8'd172 : sinpow <= 607 ;
		8'd173 : sinpow <= 612 ;
		8'd174 : sinpow <= 616 ;
		8'd175 : sinpow <= 621 ;
		8'd176 : sinpow <= 625 ;
		8'd177 : sinpow <= 630 ;
		8'd178 : sinpow <= 634 ;
		8'd179 : sinpow <= 639 ;
		8'd180 : sinpow <= 643 ;
		8'd181 : sinpow <= 648 ;
		8'd182 : sinpow <= 652 ;
		8'd183 : sinpow <= 657 ;
		8'd184 : sinpow <= 661 ;
		8'd185 : sinpow <= 666 ;
		8'd186 : sinpow <= 670 ;
		8'd187 : sinpow <= 675 ;
		8'd188 : sinpow <= 680 ;
		8'd189 : sinpow <= 684 ;
		8'd190 : sinpow <= 689 ;
		8'd191 : sinpow <= 693 ;
		8'd192 : sinpow <= 698 ;
		8'd193 : sinpow <= 703 ;
		8'd194 : sinpow <= 708 ;
		8'd195 : sinpow <= 712 ;
		8'd196 : sinpow <= 717 ;
		8'd197 : sinpow <= 722 ;
		8'd198 : sinpow <= 726 ;
		8'd199 : sinpow <= 731 ;
		8'd200 : sinpow <= 736 ;
		8'd201 : sinpow <= 741 ;
		8'd202 : sinpow <= 745 ;
		8'd203 : sinpow <= 750 ;
		8'd204 : sinpow <= 755 ;
		8'd205 : sinpow <= 760 ;
		8'd206 : sinpow <= 765 ;
		8'd207 : sinpow <= 770 ;
		8'd208 : sinpow <= 774 ;
		8'd209 : sinpow <= 779 ;
		8'd210 : sinpow <= 784 ;
		8'd211 : sinpow <= 789 ;
		8'd212 : sinpow <= 794 ;
		8'd213 : sinpow <= 799 ;
		8'd214 : sinpow <= 804 ;
		8'd215 : sinpow <= 809 ;
		8'd216 : sinpow <= 814 ;
		8'd217 : sinpow <= 819 ;
		8'd218 : sinpow <= 824 ;
		8'd219 : sinpow <= 829 ;
		8'd220 : sinpow <= 834 ;
		8'd221 : sinpow <= 839 ;
		8'd222 : sinpow <= 844 ;
		8'd223 : sinpow <= 849 ;
		8'd224 : sinpow <= 854 ;
		8'd225 : sinpow <= 859 ;
		8'd226 : sinpow <= 864 ;
		8'd227 : sinpow <= 869 ;
		8'd228 : sinpow <= 874 ;
		8'd229 : sinpow <= 880 ;
		8'd230 : sinpow <= 885 ;
		8'd231 : sinpow <= 890 ;
		8'd232 : sinpow <= 895 ;
		8'd233 : sinpow <= 900 ;
		8'd234 : sinpow <= 906 ;
		8'd235 : sinpow <= 911 ;
		8'd236 : sinpow <= 916 ;
		8'd237 : sinpow <= 921 ;
		8'd238 : sinpow <= 927 ;
		8'd239 : sinpow <= 932 ;
		8'd240 : sinpow <= 937 ;
		8'd241 : sinpow <= 942 ;
		8'd242 : sinpow <= 948 ;
		8'd243 : sinpow <= 953 ;
		8'd244 : sinpow <= 959 ;
		8'd245 : sinpow <= 964 ;
		8'd246 : sinpow <= 969 ;
		8'd247 : sinpow <= 975 ;
		8'd248 : sinpow <= 980 ;
		8'd249 : sinpow <= 986 ;
		8'd250 : sinpow <= 991 ;
		8'd251 : sinpow <= 996 ;
		8'd252 : sinpow <= 1002 ;
		8'd253 : sinpow <= 1007 ;
		8'd254 : sinpow <= 1013 ;
		8'd255 : sinpow <= 1018 ;

	endcase
end


endmodule
