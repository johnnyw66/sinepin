module musicROM  (
	input clk,
	input [8:0] address,
	output reg [7:0] note
);

always @(posedge clk)
case(address[8:0])
	  0: note<= 8'd61;
	  1: note<= 8'd63;
	  2: note<= 8'd63;
	  3: note<= 8'd61;
	  4: note<= 8'd58;
	  5: note<= 8'd58;
	  6: note<= 8'd66;
	  7: note<= 8'd66;
	  8: note<= 8'd63;
	  9: note<= 8'd63;
	 10: note<= 8'd61;
	 11: note<= 8'd61;
	 12: note<= 8'd61;
	 13: note<= 8'd61;
	 14: note<= 8'd61;
	 15: note<= 8'd61;
	 16: note<= 8'd61;
	 17: note<= 8'd63;
	 18: note<= 8'd61;
	 19: note<= 8'd63;
	 20: note<= 8'd61;
	 21: note<= 8'd61;
	 22: note<= 8'd66;
	 23: note<= 8'd66;
	 24: note<= 8'd65;
	 25: note<= 8'd65;
	 26: note<= 8'd65;
	 27: note<= 8'd65;
	 28: note<= 8'd65;
	 29: note<= 8'd65;
	 30: note<= 8'd65;
	 31: note<= 8'd65;
	 32: note<= 8'd59;
	 33: note<= 8'd61;
	 34: note<= 8'd61;
	 35: note<= 8'd59;
	 36: note<= 8'd56;
	 37: note<= 8'd56;
	 38: note<= 8'd65;
	 39: note<= 8'd65;
	 40: note<= 8'd63;
	 41: note<= 8'd63;
	 42: note<= 8'd61;
	 43: note<= 8'd61;
	 44: note<= 8'd61;
	 45: note<= 8'd61;
	 46: note<= 8'd61;
	 47: note<= 8'd61;
	 48: note<= 8'd61;
	 49: note<= 8'd63;
	 50: note<= 8'd61;
	 51: note<= 8'd63;
	 52: note<= 8'd61;
	 53: note<= 8'd61;
	 54: note<= 8'd63;
	 55: note<= 8'd63;
	 56: note<= 8'd58;
	 57: note<= 8'd58;
	 58: note<= 8'd58;
	 59: note<= 8'd58;
	 60: note<= 8'd58;
	 61: note<= 8'd58;
	 62: note<= 8'd58;
	 63: note<= 8'd58;
	 64: note<= 8'd61;
	 65: note<= 8'd63;
	 66: note<= 8'd63;
	 67: note<= 8'd61;
	 68: note<= 8'd58;
	 69: note<= 8'd58;
	 70: note<= 8'd66;
	 71: note<= 8'd66;
	 72: note<= 8'd63;
	 73: note<= 8'd63;
	 74: note<= 8'd61;
	 75: note<= 8'd61;
	 76: note<= 8'd61;
	 77: note<= 8'd61;
	 78: note<= 8'd61;
	 79: note<= 8'd61;
	 80: note<= 8'd61;
	 81: note<= 8'd63;
	 82: note<= 8'd61;
	 83: note<= 8'd63;
	 84: note<= 8'd61;
	 85: note<= 8'd61;
	 86: note<= 8'd66;
	 87: note<= 8'd66;
	 88: note<= 8'd65;
	 89: note<= 8'd65;
	 90: note<= 8'd65;
	 91: note<= 8'd65;
	 92: note<= 8'd65;
	 93: note<= 8'd65;
	 94: note<= 8'd65;
	 95: note<= 8'd65;
	 96: note<= 8'd59;
	 97: note<= 8'd61;
	 98: note<= 8'd61;
	 99: note<= 8'd59;
	100: note<= 8'd56;
	101: note<= 8'd56;
	102: note<= 8'd65;
	103: note<= 8'd65;
	104: note<= 8'd63;
	105: note<= 8'd63;
	106: note<= 8'd61;
	107: note<= 8'd61;
	108: note<= 8'd61;
	109: note<= 8'd61;
	110: note<= 8'd61;
	111: note<= 8'd61;
	112: note<= 8'd61;
	113: note<= 8'd63;
	114: note<= 8'd61;
	115: note<= 8'd63;
	116: note<= 8'd61;
	117: note<= 8'd61;
	118: note<= 8'd68;
	119: note<= 8'd68;
	120: note<= 8'd66;
	121: note<= 8'd66;
	122: note<= 8'd66;
	123: note<= 8'd66;
	124: note<= 8'd66;
	125: note<= 8'd66;
	126: note<= 8'd66;
	127: note<= 8'd66;
	128: note<= 8'd63;
	129: note<= 8'd63;
	130: note<= 8'd63;
	131: note<= 8'd63;
	132: note<= 8'd66;
	133: note<= 8'd66;
	134: note<= 8'd66;
	135: note<= 8'd63;
	136: note<= 8'd61;
	137: note<= 8'd61;
	138: note<= 8'd58;
	139: note<= 8'd58;
	140: note<= 8'd61;
	141: note<= 8'd61;
	142: note<= 8'd61;
	143: note<= 8'd61;
	144: note<= 8'd59;
	145: note<= 8'd59;
	146: note<= 8'd63;
	147: note<= 8'd63;
	148: note<= 8'd61;
	149: note<= 8'd61;
	150: note<= 8'd59;
	151: note<= 8'd59;
	152: note<= 8'd58;
	153: note<= 8'd58;
	154: note<= 8'd58;
	155: note<= 8'd58;
	156: note<= 8'd58;
	157: note<= 8'd58;
	158: note<= 8'd58;
	159: note<= 8'd58;
	160: note<= 8'd56;
	161: note<= 8'd56;
	162: note<= 8'd58;
	163: note<= 8'd58;
	164: note<= 8'd61;
	165: note<= 8'd61;
	166: note<= 8'd63;
	167: note<= 8'd63;
	168: note<= 8'd65;
	169: note<= 8'd65;
	170: note<= 8'd65;
	171: note<= 8'd65;
	172: note<= 8'd65;
	173: note<= 8'd65;
	174: note<= 8'd65;
	175: note<= 8'd65;
	176: note<= 8'd66;
	177: note<= 8'd66;
	178: note<= 8'd66;
	179: note<= 8'd66;
	180: note<= 8'd65;
	181: note<= 8'd65;
	182: note<= 8'd63;
	183: note<= 8'd63;
	184: note<= 8'd61;
	185: note<= 8'd61;
	186: note<= 8'd59;
	187: note<= 8'd56;
	188: note<= 8'd56;
	189: note<= 8'd56;
	190: note<= 8'd56;
	191: note<= 8'd56;
	192: note<= 8'd61;
	193: note<= 8'd63;
	194: note<= 8'd63;
	195: note<= 8'd61;
	196: note<= 8'd58;
	197: note<= 8'd58;
	198: note<= 8'd66;
	199: note<= 8'd66;
	200: note<= 8'd63;
	201: note<= 8'd63;
	202: note<= 8'd61;
	203: note<= 8'd61;
	204: note<= 8'd61;
	205: note<= 8'd61;
	206: note<= 8'd61;
	207: note<= 8'd61;
	208: note<= 8'd61;
	209: note<= 8'd63;
	210: note<= 8'd61;
	211: note<= 8'd63;
	212: note<= 8'd61;
	213: note<= 8'd61;
	214: note<= 8'd66;
	215: note<= 8'd66;
	216: note<= 8'd65;
	217: note<= 8'd65;
	218: note<= 8'd65;
	219: note<= 8'd65;
	220: note<= 8'd65;
	221: note<= 8'd65;
	222: note<= 8'd65;
	223: note<= 8'd65;
	224: note<= 8'd59;
	225: note<= 8'd61;
	226: note<= 8'd61;
	227: note<= 8'd59;
	228: note<= 8'd56;
	229: note<= 8'd56;
	230: note<= 8'd65;
	231: note<= 8'd65;
	232: note<= 8'd63;
	233: note<= 8'd63;
	234: note<= 8'd61;
	235: note<= 8'd61;
	236: note<= 8'd61;
	237: note<= 8'd61;
	238: note<= 8'd61;
	239: note<= 8'd61;
	240: note<= 8'd61;
	241: note<= 8'd1;
	242: note<= 8'd1;
	243: note<= 8'd1;
	244: note<= 8'd1;
	245: note<= 8'd1;
	246: note<= 8'd1;
	247: note<= 8'd1;
	248: note<= 8'd1;
	249: note<= 8'd1;
	250: note<= 8'd1;
	default: note <= 8'd0;
endcase
endmodule
