module sineCosROM #(parameter SINEROMSIZE = 256)(
	input clk,
	input [$clog2(SINEROMSIZE) - 1:0] address,
	output reg [15:0] svalue
);

always @(posedge clk)
begin
	case(address)
			8'd0 : svalue <= 16'd32768 ;
			8'd1 : svalue <= 16'd35179 ;
			8'd2 : svalue <= 16'd37523 ;
			8'd3 : svalue <= 16'd39735 ;
			8'd4 : svalue <= 16'd41753 ;
			8'd5 : svalue <= 16'd43521 ;
			8'd6 : svalue <= 16'd44988 ;
			8'd7 : svalue <= 16'd46112 ;
			8'd8 : svalue <= 16'd46857 ;
			8'd9 : svalue <= 16'd47202 ;
			8'd10 : svalue <= 16'd47130 ;
			8'd11 : svalue <= 16'd46640 ;
			8'd12 : svalue <= 16'd45738 ;
			8'd13 : svalue <= 16'd44443 ;
			8'd14 : svalue <= 16'd42783 ;
			8'd15 : svalue <= 16'd40795 ;
			8'd16 : svalue <= 16'd38524 ;
			8'd17 : svalue <= 16'd36025 ;
			8'd18 : svalue <= 16'd33356 ;
			8'd19 : svalue <= 16'd30579 ;
			8'd20 : svalue <= 16'd27763 ;
			8'd21 : svalue <= 16'd24972 ;
			8'd22 : svalue <= 16'd22275 ;
			8'd23 : svalue <= 16'd19734 ;
			8'd24 : svalue <= 16'd17410 ;
			8'd25 : svalue <= 16'd15359 ;
			8'd26 : svalue <= 16'd13626 ;
			8'd27 : svalue <= 16'd12252 ;
			8'd28 : svalue <= 16'd11267 ;
			8'd29 : svalue <= 16'd10691 ;
			8'd30 : svalue <= 16'd10535 ;
			8'd31 : svalue <= 16'd10797 ;
			8'd32 : svalue <= 16'd11466 ;
			8'd33 : svalue <= 16'd12520 ;
			8'd34 : svalue <= 16'd13928 ;
			8'd35 : svalue <= 16'd15648 ;
			8'd36 : svalue <= 16'd17632 ;
			8'd37 : svalue <= 16'd19825 ;
			8'd38 : svalue <= 16'd22166 ;
			8'd39 : svalue <= 16'd24589 ;
			8'd40 : svalue <= 16'd27030 ;
			8'd41 : svalue <= 16'd29420 ;
			8'd42 : svalue <= 16'd31694 ;
			8'd43 : svalue <= 16'd33789 ;
			8'd44 : svalue <= 16'd35647 ;
			8'd45 : svalue <= 16'd37217 ;
			8'd46 : svalue <= 16'd38453 ;
			8'd47 : svalue <= 16'd39320 ;
			8'd48 : svalue <= 16'd39792 ;
			8'd49 : svalue <= 16'd39850 ;
			8'd50 : svalue <= 16'd39491 ;
			8'd51 : svalue <= 16'd38719 ;
			8'd52 : svalue <= 16'd37550 ;
			8'd53 : svalue <= 16'd36009 ;
			8'd54 : svalue <= 16'd34132 ;
			8'd55 : svalue <= 16'd31962 ;
			8'd56 : svalue <= 16'd29552 ;
			8'd57 : svalue <= 16'd26959 ;
			8'd58 : svalue <= 16'd24245 ;
			8'd59 : svalue <= 16'd21476 ;
			8'd60 : svalue <= 16'd18719 ;
			8'd61 : svalue <= 16'd16041 ;
			8'd62 : svalue <= 16'd13506 ;
			8'd63 : svalue <= 16'd11176 ;
			8'd64 : svalue <= 16'd9107 ;
			8'd65 : svalue <= 16'd7347 ;
			8'd66 : svalue <= 16'd5939 ;
			8'd67 : svalue <= 16'd4915 ;
			8'd68 : svalue <= 16'd4298 ;
			8'd69 : svalue <= 16'd4099 ;
			8'd70 : svalue <= 16'd4321 ;
			8'd71 : svalue <= 16'd4954 ;
			8'd72 : svalue <= 16'd5980 ;
			8'd73 : svalue <= 16'd7368 ;
			8'd74 : svalue <= 16'd9079 ;
			8'd75 : svalue <= 16'd11068 ;
			8'd76 : svalue <= 16'd13279 ;
			8'd77 : svalue <= 16'd15653 ;
			8'd78 : svalue <= 16'd18127 ;
			8'd79 : svalue <= 16'd20633 ;
			8'd80 : svalue <= 16'd23106 ;
			8'd81 : svalue <= 16'd25478 ;
			8'd82 : svalue <= 16'd27687 ;
			8'd83 : svalue <= 16'd29673 ;
			8'd84 : svalue <= 16'd31381 ;
			8'd85 : svalue <= 16'd32767 ;
			8'd86 : svalue <= 16'd33792 ;
			8'd87 : svalue <= 16'd34428 ;
			8'd88 : svalue <= 16'd34654 ;
			8'd89 : svalue <= 16'd34464 ;
			8'd90 : svalue <= 16'd33860 ;
			8'd91 : svalue <= 16'd32854 ;
			8'd92 : svalue <= 16'd31471 ;
			8'd93 : svalue <= 16'd29743 ;
			8'd94 : svalue <= 16'd27713 ;
			8'd95 : svalue <= 16'd25431 ;
			8'd96 : svalue <= 16'd22952 ;
			8'd97 : svalue <= 16'd20339 ;
			8'd98 : svalue <= 16'd17656 ;
			8'd99 : svalue <= 16'd14970 ;
			8'd100 : svalue <= 16'd12348 ;
			8'd101 : svalue <= 16'd9856 ;
			8'd102 : svalue <= 16'd7555 ;
			8'd103 : svalue <= 16'd5503 ;
			8'd104 : svalue <= 16'd3751 ;
			8'd105 : svalue <= 16'd2343 ;
			8'd106 : svalue <= 16'd1312 ;
			8'd107 : svalue <= 16'd683 ;
			8'd108 : svalue <= 16'd473 ;
			8'd109 : svalue <= 16'd684 ;
			8'd110 : svalue <= 16'd1310 ;
			8'd111 : svalue <= 16'd2334 ;
			8'd112 : svalue <= 16'd3729 ;
			8'd113 : svalue <= 16'd5458 ;
			8'd114 : svalue <= 16'd7476 ;
			8'd115 : svalue <= 16'd9730 ;
			8'd116 : svalue <= 16'd12161 ;
			8'd117 : svalue <= 16'd14707 ;
			8'd118 : svalue <= 16'd17303 ;
			8'd119 : svalue <= 16'd19880 ;
			8'd120 : svalue <= 16'd22372 ;
			8'd121 : svalue <= 16'd24715 ;
			8'd122 : svalue <= 16'd26849 ;
			8'd123 : svalue <= 16'd28718 ;
			8'd124 : svalue <= 16'd30275 ;
			8'd125 : svalue <= 16'd31479 ;
			8'd126 : svalue <= 16'd32300 ;
			8'd127 : svalue <= 16'd32715 ;
			8'd128 : svalue <= 16'd32715 ;
			8'd129 : svalue <= 16'd32300 ;
			8'd130 : svalue <= 16'd31479 ;
			8'd131 : svalue <= 16'd30275 ;
			8'd132 : svalue <= 16'd28718 ;
			8'd133 : svalue <= 16'd26849 ;
			8'd134 : svalue <= 16'd24715 ;
			8'd135 : svalue <= 16'd22372 ;
			8'd136 : svalue <= 16'd19880 ;
			8'd137 : svalue <= 16'd17303 ;
			8'd138 : svalue <= 16'd14707 ;
			8'd139 : svalue <= 16'd12161 ;
			8'd140 : svalue <= 16'd9730 ;
			8'd141 : svalue <= 16'd7476 ;
			8'd142 : svalue <= 16'd5458 ;
			8'd143 : svalue <= 16'd3729 ;
			8'd144 : svalue <= 16'd2334 ;
			8'd145 : svalue <= 16'd1310 ;
			8'd146 : svalue <= 16'd684 ;
			8'd147 : svalue <= 16'd473 ;
			8'd148 : svalue <= 16'd683 ;
			8'd149 : svalue <= 16'd1312 ;
			8'd150 : svalue <= 16'd2343 ;
			8'd151 : svalue <= 16'd3751 ;
			8'd152 : svalue <= 16'd5503 ;
			8'd153 : svalue <= 16'd7555 ;
			8'd154 : svalue <= 16'd9856 ;
			8'd155 : svalue <= 16'd12348 ;
			8'd156 : svalue <= 16'd14970 ;
			8'd157 : svalue <= 16'd17656 ;
			8'd158 : svalue <= 16'd20339 ;
			8'd159 : svalue <= 16'd22952 ;
			8'd160 : svalue <= 16'd25431 ;
			8'd161 : svalue <= 16'd27713 ;
			8'd162 : svalue <= 16'd29743 ;
			8'd163 : svalue <= 16'd31471 ;
			8'd164 : svalue <= 16'd32854 ;
			8'd165 : svalue <= 16'd33860 ;
			8'd166 : svalue <= 16'd34464 ;
			8'd167 : svalue <= 16'd34654 ;
			8'd168 : svalue <= 16'd34428 ;
			8'd169 : svalue <= 16'd33792 ;
			8'd170 : svalue <= 16'd32768 ;
			8'd171 : svalue <= 16'd31381 ;
			8'd172 : svalue <= 16'd29673 ;
			8'd173 : svalue <= 16'd27687 ;
			8'd174 : svalue <= 16'd25478 ;
			8'd175 : svalue <= 16'd23106 ;
			8'd176 : svalue <= 16'd20633 ;
			8'd177 : svalue <= 16'd18127 ;
			8'd178 : svalue <= 16'd15653 ;
			8'd179 : svalue <= 16'd13279 ;
			8'd180 : svalue <= 16'd11068 ;
			8'd181 : svalue <= 16'd9079 ;
			8'd182 : svalue <= 16'd7368 ;
			8'd183 : svalue <= 16'd5980 ;
			8'd184 : svalue <= 16'd4954 ;
			8'd185 : svalue <= 16'd4321 ;
			8'd186 : svalue <= 16'd4099 ;
			8'd187 : svalue <= 16'd4298 ;
			8'd188 : svalue <= 16'd4915 ;
			8'd189 : svalue <= 16'd5939 ;
			8'd190 : svalue <= 16'd7347 ;
			8'd191 : svalue <= 16'd9107 ;
			8'd192 : svalue <= 16'd11176 ;
			8'd193 : svalue <= 16'd13506 ;
			8'd194 : svalue <= 16'd16041 ;
			8'd195 : svalue <= 16'd18719 ;
			8'd196 : svalue <= 16'd21476 ;
			8'd197 : svalue <= 16'd24245 ;
			8'd198 : svalue <= 16'd26959 ;
			8'd199 : svalue <= 16'd29552 ;
			8'd200 : svalue <= 16'd31962 ;
			8'd201 : svalue <= 16'd34132 ;
			8'd202 : svalue <= 16'd36009 ;
			8'd203 : svalue <= 16'd37550 ;
			8'd204 : svalue <= 16'd38719 ;
			8'd205 : svalue <= 16'd39491 ;
			8'd206 : svalue <= 16'd39850 ;
			8'd207 : svalue <= 16'd39792 ;
			8'd208 : svalue <= 16'd39320 ;
			8'd209 : svalue <= 16'd38453 ;
			8'd210 : svalue <= 16'd37217 ;
			8'd211 : svalue <= 16'd35647 ;
			8'd212 : svalue <= 16'd33789 ;
			8'd213 : svalue <= 16'd31694 ;
			8'd214 : svalue <= 16'd29420 ;
			8'd215 : svalue <= 16'd27030 ;
			8'd216 : svalue <= 16'd24589 ;
			8'd217 : svalue <= 16'd22166 ;
			8'd218 : svalue <= 16'd19825 ;
			8'd219 : svalue <= 16'd17632 ;
			8'd220 : svalue <= 16'd15648 ;
			8'd221 : svalue <= 16'd13928 ;
			8'd222 : svalue <= 16'd12520 ;
			8'd223 : svalue <= 16'd11466 ;
			8'd224 : svalue <= 16'd10797 ;
			8'd225 : svalue <= 16'd10535 ;
			8'd226 : svalue <= 16'd10691 ;
			8'd227 : svalue <= 16'd11267 ;
			8'd228 : svalue <= 16'd12252 ;
			8'd229 : svalue <= 16'd13626 ;
			8'd230 : svalue <= 16'd15359 ;
			8'd231 : svalue <= 16'd17410 ;
			8'd232 : svalue <= 16'd19734 ;
			8'd233 : svalue <= 16'd22275 ;
			8'd234 : svalue <= 16'd24972 ;
			8'd235 : svalue <= 16'd27763 ;
			8'd236 : svalue <= 16'd30579 ;
			8'd237 : svalue <= 16'd33356 ;
			8'd238 : svalue <= 16'd36025 ;
			8'd239 : svalue <= 16'd38524 ;
			8'd240 : svalue <= 16'd40795 ;
			8'd241 : svalue <= 16'd42783 ;
			8'd242 : svalue <= 16'd44443 ;
			8'd243 : svalue <= 16'd45738 ;
			8'd244 : svalue <= 16'd46640 ;
			8'd245 : svalue <= 16'd47130 ;
			8'd246 : svalue <= 16'd47202 ;
			8'd247 : svalue <= 16'd46857 ;
			8'd248 : svalue <= 16'd46112 ;
			8'd249 : svalue <= 16'd44988 ;
			8'd250 : svalue <= 16'd43521 ;
			8'd251 : svalue <= 16'd41753 ;
			8'd252 : svalue <= 16'd39735 ;
			8'd253 : svalue <= 16'd37523 ;
			8'd254 : svalue <= 16'd35179 ;
			8'd255 : svalue <= 16'd32768 ;
	
	endcase
end
endmodule
