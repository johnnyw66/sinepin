// SineROM case statement was generated using a simple
// bit of python
// Rather wasteful - since we only really need to produce a 
// a quarter wave of the 1st quadrant of a sine wave
// The remaining 3 quadrants are (a) reflection(s) of the 1st quadrant!

// Note: If you do make quarter sine wave tables - change
// the inapproriately named 'SINEROMSIZE' parameter - which
// is infact the number of steps taken to complete a full sinewave.
// For this particular 'ROM' - our ROM size of 256 is a complete cycle
// i.e SINEROMSIZE = 'size of ROM' = number of steps to complete a full wave.
// 'SINEROMSIZE' is the number of steps we make to complete a full wave.

/*

import math ;

fpmult = 65536 ;		#16bit
for i in range (256):
    a = i ;	
    sv = 0.5 * ( 1 + math.sin(2 * a * math.pi / 255)) ;
    fpsv =  int(fpmult * sv) ;
    # print("%d %d %d" % (i,fpsv, int(fpsv / 256))) ;
    print("8'd%d : svalue <= 16'd%d ;" % (i,fpsv)) ;

*/

module sineROM #(parameter SINEROMSIZE = 256)(
	input clk,
	input [$clog2(SINEROMSIZE) - 1:0] address,
	output  reg [15:0] svalue
);


always @(posedge clk)
begin
	case(address)

		8'd0 : svalue <= 16'd32768 ;
		8'd1 : svalue <= 16'd33575 ;
		8'd2 : svalue <= 16'd34382 ;
		8'd3 : svalue <= 16'd35187 ;
		8'd4 : svalue <= 16'd35992 ;
		8'd5 : svalue <= 16'd36794 ;
		8'd6 : svalue <= 16'd37594 ;
		8'd7 : svalue <= 16'd38391 ;
		8'd8 : svalue <= 16'd39185 ;
		8'd9 : svalue <= 16'd39975 ;
		8'd10 : svalue <= 16'd40760 ;
		8'd11 : svalue <= 16'd41541 ;
		8'd12 : svalue <= 16'd42316 ;
		8'd13 : svalue <= 16'd43085 ;
		8'd14 : svalue <= 16'd43848 ;
		8'd15 : svalue <= 16'd44605 ;
		8'd16 : svalue <= 16'd45354 ;
		8'd17 : svalue <= 16'd46095 ;
		8'd18 : svalue <= 16'd46829 ;
		8'd19 : svalue <= 16'd47554 ;
		8'd20 : svalue <= 16'd48270 ;
		8'd21 : svalue <= 16'd48976 ;
		8'd22 : svalue <= 16'd49673 ;
		8'd23 : svalue <= 16'd50360 ;
		8'd24 : svalue <= 16'd51035 ;
		8'd25 : svalue <= 16'd51700 ;
		8'd26 : svalue <= 16'd52353 ;
		8'd27 : svalue <= 16'd52994 ;
		8'd28 : svalue <= 16'd53623 ;
		8'd29 : svalue <= 16'd54240 ;
		8'd30 : svalue <= 16'd54843 ;
		8'd31 : svalue <= 16'd55433 ;
		8'd32 : svalue <= 16'd56009 ;
		8'd33 : svalue <= 16'd56571 ;
		8'd34 : svalue <= 16'd57119 ;
		8'd35 : svalue <= 16'd57652 ;
		8'd36 : svalue <= 16'd58169 ;
		8'd37 : svalue <= 16'd58672 ;
		8'd38 : svalue <= 16'd59158 ;
		8'd39 : svalue <= 16'd59629 ;
		8'd40 : svalue <= 16'd60083 ;
		8'd41 : svalue <= 16'd60521 ;
		8'd42 : svalue <= 16'd60941 ;
		8'd43 : svalue <= 16'd61345 ;
		8'd44 : svalue <= 16'd61731 ;
		8'd45 : svalue <= 16'd62100 ;
		8'd46 : svalue <= 16'd62451 ;
		8'd47 : svalue <= 16'd62784 ;
		8'd48 : svalue <= 16'd63099 ;
		8'd49 : svalue <= 16'd63395 ;
		8'd50 : svalue <= 16'd63673 ;
		8'd51 : svalue <= 16'd63932 ;
		8'd52 : svalue <= 16'd64172 ;
		8'd53 : svalue <= 16'd64393 ;
		8'd54 : svalue <= 16'd64594 ;
		8'd55 : svalue <= 16'd64777 ;
		8'd56 : svalue <= 16'd64940 ;
		8'd57 : svalue <= 16'd65083 ;
		8'd58 : svalue <= 16'd65207 ;
		8'd59 : svalue <= 16'd65311 ;
		8'd60 : svalue <= 16'd65396 ;
		8'd61 : svalue <= 16'd65460 ;
		8'd62 : svalue <= 16'd65505 ;
		8'd63 : svalue <= 16'd65530 ;
		8'd64 : svalue <= 16'd65535 ;
		8'd65 : svalue <= 16'd65520 ;
		8'd66 : svalue <= 16'd65485 ;
		8'd67 : svalue <= 16'd65430 ;
		8'd68 : svalue <= 16'd65356 ;
		8'd69 : svalue <= 16'd65262 ;
		8'd70 : svalue <= 16'd65148 ;
		8'd71 : svalue <= 16'd65014 ;
		8'd72 : svalue <= 16'd64861 ;
		8'd73 : svalue <= 16'd64688 ;
		8'd74 : svalue <= 16'd64496 ;
		8'd75 : svalue <= 16'd64285 ;
		8'd76 : svalue <= 16'd64054 ;
		8'd77 : svalue <= 16'd63805 ;
		8'd78 : svalue <= 16'd63536 ;
		8'd79 : svalue <= 16'd63249 ;
		8'd80 : svalue <= 16'd62944 ;
		8'd81 : svalue <= 16'd62620 ;
		8'd82 : svalue <= 16'd62278 ;
		8'd83 : svalue <= 16'd61918 ;
		8'd84 : svalue <= 16'd61540 ;
		8'd85 : svalue <= 16'd61145 ;
		8'd86 : svalue <= 16'd60733 ;
		8'd87 : svalue <= 16'd60304 ;
		8'd88 : svalue <= 16'd59858 ;
		8'd89 : svalue <= 16'd59396 ;
		8'd90 : svalue <= 16'd58917 ;
		8'd91 : svalue <= 16'd58422 ;
		8'd92 : svalue <= 16'd57912 ;
		8'd93 : svalue <= 16'd57387 ;
		8'd94 : svalue <= 16'd56847 ;
		8'd95 : svalue <= 16'd56292 ;
		8'd96 : svalue <= 16'd55723 ;
		8'd97 : svalue <= 16'd55140 ;
		8'd98 : svalue <= 16'd54543 ;
		8'd99 : svalue <= 16'd53933 ;
		8'd100 : svalue <= 16'd53311 ;
		8'd101 : svalue <= 16'd52675 ;
		8'd102 : svalue <= 16'd52028 ;
		8'd103 : svalue <= 16'd51369 ;
		8'd104 : svalue <= 16'd50699 ;
		8'd105 : svalue <= 16'd50018 ;
		8'd106 : svalue <= 16'd49326 ;
		8'd107 : svalue <= 16'd48624 ;
		8'd108 : svalue <= 16'd47913 ;
		8'd109 : svalue <= 16'd47192 ;
		8'd110 : svalue <= 16'd46463 ;
		8'd111 : svalue <= 16'd45726 ;
		8'd112 : svalue <= 16'd44980 ;
		8'd113 : svalue <= 16'd44227 ;
		8'd114 : svalue <= 16'd43468 ;
		8'd115 : svalue <= 16'd42701 ;
		8'd116 : svalue <= 16'd41929 ;
		8'd117 : svalue <= 16'd41151 ;
		8'd118 : svalue <= 16'd40368 ;
		8'd119 : svalue <= 16'd39580 ;
		8'd120 : svalue <= 16'd38789 ;
		8'd121 : svalue <= 16'd37993 ;
		8'd122 : svalue <= 16'd37195 ;
		8'd123 : svalue <= 16'd36393 ;
		8'd124 : svalue <= 16'd35590 ;
		8'd125 : svalue <= 16'd34785 ;
		8'd126 : svalue <= 16'd33978 ;
		8'd127 : svalue <= 16'd33171 ;
		8'd128 : svalue <= 16'd32364 ;
		8'd129 : svalue <= 16'd31557 ;
		8'd130 : svalue <= 16'd30750 ;
		8'd131 : svalue <= 16'd29945 ;
		8'd132 : svalue <= 16'd29142 ;
		8'd133 : svalue <= 16'd28340 ;
		8'd134 : svalue <= 16'd27542 ;
		8'd135 : svalue <= 16'd26746 ;
		8'd136 : svalue <= 16'd25955 ;
		8'd137 : svalue <= 16'd25167 ;
		8'd138 : svalue <= 16'd24384 ;
		8'd139 : svalue <= 16'd23606 ;
		8'd140 : svalue <= 16'd22834 ;
		8'd141 : svalue <= 16'd22067 ;
		8'd142 : svalue <= 16'd21308 ;
		8'd143 : svalue <= 16'd20555 ;
		8'd144 : svalue <= 16'd19809 ;
		8'd145 : svalue <= 16'd19072 ;
		8'd146 : svalue <= 16'd18343 ;
		8'd147 : svalue <= 16'd17622 ;
		8'd148 : svalue <= 16'd16911 ;
		8'd149 : svalue <= 16'd16209 ;
		8'd150 : svalue <= 16'd15517 ;
		8'd151 : svalue <= 16'd14836 ;
		8'd152 : svalue <= 16'd14166 ;
		8'd153 : svalue <= 16'd13507 ;
		8'd154 : svalue <= 16'd12860 ;
		8'd155 : svalue <= 16'd12224 ;
		8'd156 : svalue <= 16'd11602 ;
		8'd157 : svalue <= 16'd10992 ;
		8'd158 : svalue <= 16'd10395 ;
		8'd159 : svalue <= 16'd9812 ;
		8'd160 : svalue <= 16'd9243 ;
		8'd161 : svalue <= 16'd8688 ;
		8'd162 : svalue <= 16'd8148 ;
		8'd163 : svalue <= 16'd7623 ;
		8'd164 : svalue <= 16'd7113 ;
		8'd165 : svalue <= 16'd6618 ;
		8'd166 : svalue <= 16'd6139 ;
		8'd167 : svalue <= 16'd5677 ;
		8'd168 : svalue <= 16'd5231 ;
		8'd169 : svalue <= 16'd4802 ;
		8'd170 : svalue <= 16'd4390 ;
		8'd171 : svalue <= 16'd3995 ;
		8'd172 : svalue <= 16'd3617 ;
		8'd173 : svalue <= 16'd3257 ;
		8'd174 : svalue <= 16'd2915 ;
		8'd175 : svalue <= 16'd2591 ;
		8'd176 : svalue <= 16'd2286 ;
		8'd177 : svalue <= 16'd1999 ;
		8'd178 : svalue <= 16'd1730 ;
		8'd179 : svalue <= 16'd1481 ;
		8'd180 : svalue <= 16'd1250 ;
		8'd181 : svalue <= 16'd1039 ;
		8'd182 : svalue <= 16'd847 ;
		8'd183 : svalue <= 16'd674 ;
		8'd184 : svalue <= 16'd521 ;
		8'd185 : svalue <= 16'd387 ;
		8'd186 : svalue <= 16'd273 ;
		8'd187 : svalue <= 16'd179 ;
		8'd188 : svalue <= 16'd105 ;
		8'd189 : svalue <= 16'd50 ;
		8'd190 : svalue <= 16'd15 ;
		8'd191 : svalue <= 16'd0 ;
		8'd192 : svalue <= 16'd5 ;
		8'd193 : svalue <= 16'd30 ;
		8'd194 : svalue <= 16'd75 ;
		8'd195 : svalue <= 16'd139 ;
		8'd196 : svalue <= 16'd224 ;
		8'd197 : svalue <= 16'd328 ;
		8'd198 : svalue <= 16'd452 ;
		8'd199 : svalue <= 16'd595 ;
		8'd200 : svalue <= 16'd758 ;
		8'd201 : svalue <= 16'd941 ;
		8'd202 : svalue <= 16'd1142 ;
		8'd203 : svalue <= 16'd1363 ;
		8'd204 : svalue <= 16'd1603 ;
		8'd205 : svalue <= 16'd1862 ;
		8'd206 : svalue <= 16'd2140 ;
		8'd207 : svalue <= 16'd2436 ;
		8'd208 : svalue <= 16'd2751 ;
		8'd209 : svalue <= 16'd3084 ;
		8'd210 : svalue <= 16'd3435 ;
		8'd211 : svalue <= 16'd3804 ;
		8'd212 : svalue <= 16'd4190 ;
		8'd213 : svalue <= 16'd4594 ;
		8'd214 : svalue <= 16'd5014 ;
		8'd215 : svalue <= 16'd5452 ;
		8'd216 : svalue <= 16'd5906 ;
		8'd217 : svalue <= 16'd6377 ;
		8'd218 : svalue <= 16'd6863 ;
		8'd219 : svalue <= 16'd7366 ;
		8'd220 : svalue <= 16'd7883 ;
		8'd221 : svalue <= 16'd8416 ;
		8'd222 : svalue <= 16'd8964 ;
		8'd223 : svalue <= 16'd9526 ;
		8'd224 : svalue <= 16'd10102 ;
		8'd225 : svalue <= 16'd10692 ;
		8'd226 : svalue <= 16'd11295 ;
		8'd227 : svalue <= 16'd11912 ;
		8'd228 : svalue <= 16'd12541 ;
		8'd229 : svalue <= 16'd13182 ;
		8'd230 : svalue <= 16'd13835 ;
		8'd231 : svalue <= 16'd14500 ;
		8'd232 : svalue <= 16'd15175 ;
		8'd233 : svalue <= 16'd15862 ;
		8'd234 : svalue <= 16'd16559 ;
		8'd235 : svalue <= 16'd17265 ;
		8'd236 : svalue <= 16'd17981 ;
		8'd237 : svalue <= 16'd18706 ;
		8'd238 : svalue <= 16'd19440 ;
		8'd239 : svalue <= 16'd20181 ;
		8'd240 : svalue <= 16'd20930 ;
		8'd241 : svalue <= 16'd21687 ;
		8'd242 : svalue <= 16'd22450 ;
		8'd243 : svalue <= 16'd23219 ;
		8'd244 : svalue <= 16'd23994 ;
		8'd245 : svalue <= 16'd24775 ;
		8'd246 : svalue <= 16'd25560 ;
		8'd247 : svalue <= 16'd26350 ;
		8'd248 : svalue <= 16'd27144 ;
		8'd249 : svalue <= 16'd27941 ;
		8'd250 : svalue <= 16'd28741 ;
		8'd251 : svalue <= 16'd29543 ;
		8'd252 : svalue <= 16'd30348 ;
		8'd253 : svalue <= 16'd31153 ;
		8'd254 : svalue <= 16'd31960 ;
		8'd255 : svalue <= 16'd32767 ;
		//default: svalue <= 0 ;
	endcase
end
endmodule
